class sseqr_ahb extends uvm_sequencer#(slv_item_ahb);

function new(string name = "sseqr_ahb",uvm_component parent);
super.new(name,parent);
endfunction

endclass