class sequence_ahb extends uvm_sequence_item;

    `uvm_object_utils(sequence_ahb);
    

endclass