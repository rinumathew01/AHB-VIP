class slv_item_ahb extends uvm_sequence_item;

    `uvm_object_utils(slv_item_ahb);
    

endclass : slv_item_ahb