class mseqr_ahb extends uvm_sequencer#(mstr_item_ahb);

function new(string name = "mseqr_ahb",uvm_component parent);
super.new(name,parent);
endfunction

endclass