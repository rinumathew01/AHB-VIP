class mstr_seq_ahb extends uvm_sequence#(mstr_item_ahb);

    `uvm_object_utils(mstr_seq_ahb);
    

endclass : mstr_seq_ahb