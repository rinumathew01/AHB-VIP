class mstr_item_ahb extends uvm_sequence_item;

    `uvm_object_utils(mstr_item_ahb);
    

endclass : mstr_item_ahb