class env_config extends uvm_config;
    `uvm_object_utils(env_config)

endclass