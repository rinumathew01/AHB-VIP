package pkg_ahb;
    `include "uvm_macros.svh"
    import uvm_pkg::*;

    `include "intf_ahb.sv"
    `include "test_ahb.sv"
    `include "env_ahb.sv"
    `include "mstr_agnt_ahb.sv"
    `include "slv_agnt_ahb.sv"
    `include "mstr_driv_ahb.sv"
    `include "slv_driv_ahb.sv"
    `include "mstr_mon_ahb.sv"
    `include "slv_mon_ahb.sv"
    `include "sequence_ahb.sv"
    `include "seq_item_ahb.sv"

endpackage