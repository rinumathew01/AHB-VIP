class seq_item_ahb extends uvm_sequence_item;

    `uvm_object_utils(seq_item_ahb);
    

endclass