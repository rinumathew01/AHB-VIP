package pkg_ahb;
    `include "uvm_macros.svh"
    import uvm_pkg::*;

    `include "mstr_item_ahb.sv"
    `include "slv_item_ahb.sv"
    `include "mstr_seq_ahb.sv"
    `include "slv_seq_ahb.sv"
    `include "magnt_config.sv"
    `include "sagnt_config.sv"
    `include "env_config.sv"
    `include "mseqr_ahb.sv"
    `include "sseqr_ahb.sv"
    `include "vseqr_ahb.sv"
    `include "mstr_driv_ahb.sv"
    `include "slv_driv_ahb.sv"
    `include "mstr_mon_ahb.sv"
    `include "slv_mon_ahb.sv"
    `include "mstr_agnt_ahb.sv"
    `include "slv_agnt_ahb.sv"
    `include "env_ahb.sv"
    `include "test_ahb.sv"


endpackage