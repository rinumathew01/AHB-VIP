class slv_seq_ahb extends uvm_sequence_item;

    `uvm_object_utils(slv_seq_ahb);
    

endclass