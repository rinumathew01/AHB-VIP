interface intf_ahb;

endinterface